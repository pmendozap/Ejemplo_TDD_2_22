`timescale 1ns / 1ps

module fsm_pulsos();
endmodule

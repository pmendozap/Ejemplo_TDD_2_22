`timescale 1ns / 1ps

module fsm_pulsos_tb;
    fsm_pulsos dut();
endmodule;